module fsm (

input clk,
input rst,
input pause,
input 10start,
input start

){
.clk(rst){
.rst{ 
}


}
