module bcd_counter
 # (paramater SIZE = 7)
(
  output [SIZE-1:0] number,
  input logic second_tick,

)
