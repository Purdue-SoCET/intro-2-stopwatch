module tb_fsm
